// Exercise 2-1-4: AND Gate
module AND_gate (
    input a,
    input b,
    output out
);
    assign out = a & b;
endmodule