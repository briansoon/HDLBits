// Exercise 3-1-1-1: Wire
module Wire (
    input in,
    output out
);
    assign out = in;
endmodule