// Exercise 3-1-1-2: GND
module GND (
    output out
);
    assign out = 1'b0;
endmodule