// Exercise 1-2: Output Zero
module zero_out (output zero);
    assign zero = 1'b0;
endmodule