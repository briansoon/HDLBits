// Exercise 2-1-8: 7458 chip
module chip_7458 (
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y
);
    // output of AND gates = input of OR gates
    wire w1, w2, w3, w4;

    // AND gates output
    assign w1 = p2c & p2d;
    assign w2 = p2a & p2b;
    assign w3 = p1a & p1b & p1c;
    assign w4 = p1d & p1e & p1f;

    // final OR gates outputs
    assign p1y = w3 | w4;
    assign p2y = w1 | w2;

endmodule