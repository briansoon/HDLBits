// Exercise 2-1-3: Inverter
module Invert (
    input in,
    output out
);
    assign out = ~in;
endmodule