// Exercise 1-1: Getting Started
module one_out (output one);
    assign one = 1'b1;
endmodule