// Exercise 2-1-1: Simple Wire
module SimpleWire (
    input in,
    output out
);
    assign out = in;
endmodule